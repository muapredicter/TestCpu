module IO(
    input wire ce,
    input wire clk,
    input wire we,
    input wire [31:0] addr,
    input wire [31:0] wtData,
    output reg [31:0] rdData
    /*IO interface*/
);
/*access IO device*/
endmodule